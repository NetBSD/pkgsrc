@comment $NetBSD: PLIST.sv,v 1.1.1.1 2009/04/26 04:01:49 taca Exp $
${TL_WEBDIR}/system/modules/backend/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/backend/languages/sv/countries.php
${TL_WEBDIR}/system/modules/backend/languages/sv/default.php
${TL_WEBDIR}/system/modules/backend/languages/sv/explain.php
${TL_WEBDIR}/system/modules/backend/languages/sv/languages.php
${TL_WEBDIR}/system/modules/backend/languages/sv/modules.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_article.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_content.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_files.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_flash.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_form.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_form_field.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_layout.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_log.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_maintenance.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_member.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_member_group.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_page.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_settings.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_style.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_style_sheet.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_task.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_undo.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_user.php
${TL_WEBDIR}/system/modules/backend/languages/sv/tl_user_group.php
${TL_WEBDIR}/system/modules/calendar/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/calendar/languages/sv/default.php
${TL_WEBDIR}/system/modules/calendar/languages/sv/modules.php
${TL_WEBDIR}/system/modules/calendar/languages/sv/tl_calendar.php
${TL_WEBDIR}/system/modules/calendar/languages/sv/tl_calendar_events.php
${TL_WEBDIR}/system/modules/calendar/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/calendar/languages/sv/tl_user.php
${TL_WEBDIR}/system/modules/calendar/languages/sv/tl_user_group.php
${TL_WEBDIR}/system/modules/comments/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/comments/languages/sv/modules.php
${TL_WEBDIR}/system/modules/comments/languages/sv/tl_comments.php
${TL_WEBDIR}/system/modules/comments/languages/sv/tl_content.php
${TL_WEBDIR}/system/modules/dfGallery/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/dfGallery/languages/sv/default.php
${TL_WEBDIR}/system/modules/dfGallery/languages/sv/modules.php
${TL_WEBDIR}/system/modules/dfGallery/languages/sv/tl_content.php
${TL_WEBDIR}/system/modules/faq/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/faq/languages/sv/default.php
${TL_WEBDIR}/system/modules/faq/languages/sv/modules.php
${TL_WEBDIR}/system/modules/faq/languages/sv/tl_faq.php
${TL_WEBDIR}/system/modules/faq/languages/sv/tl_faq_category.php
${TL_WEBDIR}/system/modules/faq/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/frontend/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/frontend/languages/sv/default.php
${TL_WEBDIR}/system/modules/frontend/languages/sv/modules.php
${TL_WEBDIR}/system/modules/listing/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/listing/languages/sv/default.php
${TL_WEBDIR}/system/modules/listing/languages/sv/modules.php
${TL_WEBDIR}/system/modules/listing/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/memberlist/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/memberlist/languages/sv/default.php
${TL_WEBDIR}/system/modules/memberlist/languages/sv/modules.php
${TL_WEBDIR}/system/modules/memberlist/languages/sv/tl_member.php
${TL_WEBDIR}/system/modules/memberlist/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/news/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/news/languages/sv/default.php
${TL_WEBDIR}/system/modules/news/languages/sv/modules.php
${TL_WEBDIR}/system/modules/news/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/news/languages/sv/tl_news.php
${TL_WEBDIR}/system/modules/news/languages/sv/tl_news_archive.php
${TL_WEBDIR}/system/modules/news/languages/sv/tl_news_comments.php
${TL_WEBDIR}/system/modules/news/languages/sv/tl_user.php
${TL_WEBDIR}/system/modules/news/languages/sv/tl_user_group.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/newsletter/languages/sv/default.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/modules.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/tl_member.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/tl_newsletter.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/tl_newsletter_channel.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/tl_newsletter_recipients.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/tl_user.php
${TL_WEBDIR}/system/modules/newsletter/languages/sv/tl_user_group.php
${TL_WEBDIR}/system/modules/registration/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/registration/languages/sv/default.php
${TL_WEBDIR}/system/modules/registration/languages/sv/modules.php
${TL_WEBDIR}/system/modules/registration/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/rep_base/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/rep_base/languages/sv/modules.php
${TL_WEBDIR}/system/modules/rep_base/languages/sv/tl_repository.php
${TL_WEBDIR}/system/modules/rep_base/languages/sv/tl_settings.php
${TL_WEBDIR}/system/modules/rep_client/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/rep_client/languages/sv/modules.php
${TL_WEBDIR}/system/modules/rep_client/languages/sv/tl_repository.php
${TL_WEBDIR}/system/modules/rep_client/languages/sv/tl_settings.php
${TL_WEBDIR}/system/modules/rss_reader/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/rss_reader/languages/sv/modules.php
${TL_WEBDIR}/system/modules/rss_reader/languages/sv/tl_module.php
${TL_WEBDIR}/system/modules/tpl_editor/languages/sv/.htaccess
${TL_WEBDIR}/system/modules/tpl_editor/languages/sv/modules.php
${TL_WEBDIR}/system/modules/tpl_editor/languages/sv/tl_templates.php
@dirrm ${TL_WEBDIR}/system/modules/tpl_editor/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/rss_reader/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/rep_client/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/rep_base/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/registration/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/newsletter/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/news/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/memberlist/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/listing/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/frontend/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/faq/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/dfGallery/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/comments/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/calendar/languages/sv
@dirrm ${TL_WEBDIR}/system/modules/backend/languages/sv
